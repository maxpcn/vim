module clk_gate_ran(
    input       clk,
    input       genp,
    input       testmodep,
    output      gclk);


endmodule
